skxja
