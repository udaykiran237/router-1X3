askbxka
